*** SPICE deck for cell Andgate{sch} from library SP20_VlsiCEP_FA17_BCE_004_016
*** Created on Sat Jun 19, 2021 17:05:35
*** Last revised on Thu Jun 24, 2021 08:37:58
*** Written on Thu Jun 24, 2021 09:14:33 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

.global gnd vdd

*** TOP LEVEL CELL: Andgate{sch}
Mnmos-4@1 net@36 B gnd gnd N L=0.6U W=3U
Mnmos-4@2 Output A net@36 gnd N L=0.6U W=3U
Mpmos-4@0 Output B vdd vdd P L=0.6U W=3U
Mpmos-4@1 Output A vdd vdd P L=0.6U W=3U

* Spice Code nodes in cell cell 'Andgate{sch}'
vdd vdd 0 DC 5
vA A  0 pulse (0 5 0 1n 1n 10n 20n)
vB B  0 pulse (0 5 0 1n 1n 10n 20n)
.trans 1n 100n
.include C:\Program Files (x86)\Electric\C5_models.txt
.END
